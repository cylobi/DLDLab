module TopModule(
    input sel,
    input [4:0] msg,
    input rst,
    input init,
    input [2:0]sw,
    input mode,
    output out
)

