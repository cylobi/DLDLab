module Resulator(input signBit, [7:0] XIn, output reg [7:0] YOut);

wire [8:0] MSB
Twos_complement tc(.a())

endmodule