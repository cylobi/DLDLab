module SineController
(
    input clk, 
    rst,
    output reg signBit, 
    phasePos, 
    [5:0] addr, 
);

reg [63:0] sine;



endmodule